module vvcatio
