module vvcatio

import vvnet
import vvpoller

fn serve() int {
}

